library ieee;
use ieee.std_logic_1164.all;
library lattice;
use lattice.all;
library machxo2;
use machxo2.all;
use packageosc00.all;


entity init00 is
port(
	clkinit: in std_logic;
	inFlaginit: in std_logic;
	codopinit: in std_logic_vector(3 downto 0);
	outAC8init: out std_logic_vector(7 downto 0);
	outAC12init: out std_logic_vector(11 downto 0);
	outFlag12init: out std_logic;
	outFlag8init: out std_logic
);
end entity;


architecture init0 of init00 is
begin

	pinit: process(clkinit)
	variable aux0: bit:='0';
	variable aux: bit:='0';
	begin
		if(clkinit' event and clkinit= '0')then
		if(codopinit="0000") then
		case inFlaginit is
			when '1' =>
				if(aux0 = '0') then
					aux:='1';
					outAC8init <= "00111100";
					outAC12init <="000011110000";
					outFlag8init<='1';
					outFlag12init<='1';
				else
					outFlag8init<='0';
					outFlag12init<='0';
				end if;
			when '0' =>
			when others => null;
			end case;
		else
			outAC8init <= (others => 'Z');
			outAC12init <= (others => 'Z');
			outFlag8init <='Z';
			outFlag12init <='Z';
			aux0:='0';
			aux:='0';
		end if;-- cod op
		end if;
	end process pinit;
end init0;