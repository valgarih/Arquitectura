/* Verilog model created from schematic mutiplicador.sch -- Dec 08, 2015 13:40 */

module mutiplicador;




endmodule // mutiplicador
